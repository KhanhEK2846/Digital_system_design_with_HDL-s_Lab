module BCD_2_LED_7_Segment (L1,L0,X);
input [6:0]X;
output reg [3:0] L1;
output reg [3:0] L0;

always@(*)
begin
if(X < 7'd10)
begin 
	L1 <= 4'b0;
	L0 <= X;
end

if(X > 7'd9 && X < 7'd20)
begin
	L1 <= 4'd1;
	L0 <=	(X == 6'd10)? 4'd0:
			(X == 6'd11)? 4'd1 : 
			(X == 6'd12)? 4'd2 :
			(X == 6'd13)? 4'd3 :
			(X == 6'd14)? 4'd4 :
			(X == 6'd15)? 4'd5 :
			(X == 6'd16)? 4'd6 :
			(X == 6'd17)? 4'd7 :
			(X == 6'd18)? 4'd8 : 4'd9;
end

if(X > 7'd19 && X < 7'd30)
begin
	L1 <= 4'd2;
	L0 <=	(X == 6'd20)? 4'd0:
			(X == 6'd21)? 4'd1 : 
			(X == 6'd22)? 4'd2 :
			(X == 6'd23)? 4'd3 :
			(X == 6'd24)? 4'd4 :
			(X == 6'd25)? 4'd5 :
			(X == 6'd26)? 4'd6 :
			(X == 6'd27)? 4'd7 :
			(X == 6'd28)? 4'd8 : 4'd9;
end

if(X > 7'd29 && X < 7'd40)
begin
	L1 <= 4'd3;
	L0 <=	(X == 6'd30)? 4'd0:
			(X == 6'd31)? 4'd1 : 
			(X == 6'd32)? 4'd2 :
			(X == 6'd33)? 4'd3 :
			(X == 6'd34)? 4'd4 :
			(X == 6'd35)? 4'd5 :
			(X == 6'd36)? 4'd6 :
			(X == 6'd37)? 4'd7 :
			(X == 6'd38)? 4'd8 : 4'd9;
end

if(X > 7'd39 && X < 7'd50)
begin
	L1 <= 4'd4;
	L0 <=	(X == 6'd40)? 4'd0:
			(X == 6'd41)? 4'd1 : 
			(X == 6'd42)? 4'd2 :
			(X == 6'd43)? 4'd3 :
			(X == 6'd44)? 4'd4 :
			(X == 6'd45)? 4'd5 :
			(X == 6'd46)? 4'd6 :
			(X == 6'd47)? 4'd7 :
			(X == 6'd48)? 4'd8 : 4'd9;
end

if(X > 7'd49 && X < 7'd60)
begin
	L1 <= 4'd5;
	L0 <=	(X == 6'd50)? 4'd0:
			(X == 6'd51)? 4'd1 : 
			(X == 6'd52)? 4'd2 :
			(X == 6'd53)? 4'd3 :
			(X == 6'd54)? 4'd4 :
			(X == 6'd55)? 4'd5 :
			(X == 6'd56)? 4'd6 :
			(X == 6'd57)? 4'd7 :
			(X == 6'd58)? 4'd8 : 4'd9;
end

if(X > 7'd59 && X < 7'd70)
begin
	L1 <= 4'd6;
	L0 <=	(X == 6'd60)? 4'd0:
			(X == 6'd61)? 4'd1 : 
			(X == 6'd62)? 4'd2 :
			(X == 6'd63)? 4'd3 :
			(X == 6'd64)? 4'd4 :
			(X == 6'd65)? 4'd5 :
			(X == 6'd66)? 4'd6 :
			(X == 6'd67)? 4'd7 :
			(X == 6'd68)? 4'd8 : 4'd9;
end

if(X > 7'd69 && X < 7'd80)
begin
	L1 <= 4'd7;
	L0 <=	(X == 6'd70)? 4'd0:
			(X == 6'd71)? 4'd1 : 
			(X == 6'd72)? 4'd2 :
			(X == 6'd73)? 4'd3 :
			(X == 6'd74)? 4'd4 :
			(X == 6'd75)? 4'd5 :
			(X == 6'd76)? 4'd6 :
			(X == 6'd77)? 4'd7 :
			(X == 6'd78)? 4'd8 : 4'd9;
end

if(X > 7'd79 && X < 7'd90)
begin
	L1 <= 4'd8;
	L0 <=	(X == 6'd80)? 4'd0:
			(X == 6'd81)? 4'd1 : 
			(X == 6'd82)? 4'd2 :
			(X == 6'd83)? 4'd3 :
			(X == 6'd84)? 4'd4 :
			(X == 6'd85)? 4'd5 :
			(X == 6'd86)? 4'd6 :
			(X == 6'd87)? 4'd7 :
			(X == 6'd88)? 4'd8 : 4'd9;
end

if(X > 7'd89 && X < 7'd100)
begin
	L1 <= 4'd9;
	L0 <=	(X == 6'd90)? 4'd0:
			(X == 6'd91)? 4'd1 : 
			(X == 6'd92)? 4'd2 :
			(X == 6'd93)? 4'd3 :
			(X == 6'd94)? 4'd4 :
			(X == 6'd95)? 4'd5 :
			(X == 6'd96)? 4'd6 :
			(X == 6'd97)? 4'd7 :
			(X == 6'd98)? 4'd8 : 4'd9;
end

end
